module dictionary(
	input [6:0] id,
	output reg [4:0] wordnum,
	output reg [74:0] word // 5 bits per alphabet, length <= 15
);


endmodule