module dictionary(
	input id,
	output reg [74:0] word // 5 bits per alphabet, length <= 15
);


endmodule